class source_agent extends uvm_agent;
	
	`uvm_component_utils(source_agent)
	
	source_agent_config src_cfg;
	
	source_monitor monh;
	source_driver drvh;
	source_sequencer sqrh;
	
	function new(string name = "source_agent", uvm_component parent);
		super.new(name,parent);
	endfunction
	
	function void build_phase(uvm_phase phase);
		super.build_phase(phase);
		if(!uvm_config_db#(source_agent_config)::get(this,"","source_agent_config",src_cfg))
				`uvm_fatal("src_agt", "cannot get source_agent_config")
		monh = source_monitor::type_id::create("monh", this);
		if(src_cfg.is_active==UVM_ACTIVE)
			begin
				drvh = source_driver::type_id::create("drvh",this);
				sqrh = source_sequencer::type_id::create("sqrh",this);
			end
	endfunction
	
	function void connect_phase(uvm_phase phase);
		if(src_cfg.is_active==UVM_ACTIVE) begin
				drvh.seq_item_port.connect(sqrh.seq_item_export);
		end
	endfunction
	
endclass
		