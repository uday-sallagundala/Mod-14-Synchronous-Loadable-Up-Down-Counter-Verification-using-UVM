class counter_reference_model extends uvm_component;
	`uvm_component_utils(counter_reference_model)
	
	function new(string name = "counter_reference_model", uvm_component parent);
		super.new(name,parent);
	endfunction
endclass
